library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity bin2bcd is
    Port (
        bin_in : in  std_logic_vector(7 downto 0); 
        bcd0   : out std_logic_vector(3 downto 0); -- Unidade
        bcd1   : out std_logic_vector(3 downto 0); -- Dezena
        bcd2   : out std_logic_vector(3 downto 0); -- Centena
        bcd3   : out std_logic_vector(3 downto 0)  -- Milhar
    );
end entity;

architecture Behavioral of bin2bcd is

    type bcd_type is array (0 to 255) of std_logic_vector(15 downto 0);
    constant bcd: bcd_type := (
        0 => "0000000000000000",
        1 => "0000000000000001",
        2 => "0000000000000010",
        3 => "0000000000000011",
        4 => "0000000000000100",
        5 => "0000000000000101",
        6 => "0000000000000110",
        7 => "0000000000000111",
        8 => "0000000000001000",
        9 => "0000000000001001",
        10 => "0000000000010000",
        11 => "0000000000010001",
        12 => "0000000000010010",
        13 => "0000000000010011",
        14 => "0000000000010100",
        15 => "0000000000010101",
        16 => "0000000000010110",
        17 => "0000000000010111",
        18 => "0000000000011000",
        19 => "0000000000011001",
        20 => "0000000000100000",
        21 => "0000000000100001",
        22 => "0000000000100010",
        23 => "0000000000100011",
        24 => "0000000000100100",
        25 => "0000000000100101",
        26 => "0000000000100110",
        27 => "0000000000100111",
        28 => "0000000000101000",
        29 => "0000000000101001",
        30 => "0000000000110000",
        31 => "0000000000110001",
        32 => "0000000000110010",
        33 => "0000000000110011",
        34 => "0000000000110100",
        35 => "0000000000110101",
        36 => "0000000000110110",
        37 => "0000000000110111",
        38 => "0000000000111000",
        39 => "0000000000111001",
        40 => "0000000001000000",
        41 => "0000000001000001",
        42 => "0000000001000010",
        43 => "0000000001000011",
        44 => "0000000001000100",
        45 => "0000000001000101",
        46 => "0000000001000110",
        47 => "0000000001000111",
        48 => "0000000001001000",
        49 => "0000000001001001",
        50 => "0000000001010000",
        51 => "0000000001010001",
        52 => "0000000001010010",
        53 => "0000000001010011",
        54 => "0000000001010100",
        55 => "0000000001010101",
        56 => "0000000001010110",
        57 => "0000000001010111",
        58 => "0000000001011000",
        59 => "0000000001011001",
        60 => "0000000001100000",
        61 => "0000000001100001",
        62 => "0000000001100010",
        63 => "0000000001100011",
        64 => "0000000001100100",
        65 => "0000000001100101",
        66 => "0000000001100110",
        67 => "0000000001100111",
        68 => "0000000001101000",
        69 => "0000000001101001",
        70 => "0000000001110000",
        71 => "0000000001110001",
        72 => "0000000001110010",
        73 => "0000000001110011",
        74 => "0000000001110100",
        75 => "0000000001110101",
        76 => "0000000001110110",
        77 => "0000000001110111",
        78 => "0000000001111000",
        79 => "0000000001111001",
        80 => "0000000010000000",
        81 => "0000000010000001",
        82 => "0000000010000010",
        83 => "0000000010000011",
        84 => "0000000010000100",
        85 => "0000000010000101",
        86 => "0000000010000110",
        87 => "0000000010000111",
        88 => "0000000010001000",
        89 => "0000000010001001",
        90 => "0000000010010000",
        91 => "0000000010010001",
        92 => "0000000010010010",
        93 => "0000000010010011",
        94 => "0000000010010100",
        95 => "0000000010010101",
        96 => "0000000010010110",
        97 => "0000000010010111",
        98 => "0000000010011000",
        99 => "0000000010011001",
        100 => "0000000100000000",
        101 => "0000000100000001",
        102 => "0000000100000010",
        103 => "0000000100000011",
        104 => "0000000100000100",
        105 => "0000000100000101",
        106 => "0000000100000110",
        107 => "0000000100000111",
        108 => "0000000100001000",
        109 => "0000000100001001",
        110 => "0000000100010000",
        111 => "0000000100010001",
        112 => "0000000100010010",
        113 => "0000000100010011",
        114 => "0000000100010100",
        115 => "0000000100010101",
        116 => "0000000100010110",
        117 => "0000000100010111",
        118 => "0000000100011000",
        119 => "0000000100011001",
        120 => "0000000100100000",
        121 => "0000000100100001",
        122 => "0000000100100010",
        123 => "0000000100100011",
        124 => "0000000100100100",
        125 => "0000000100100101",
        126 => "0000000100100110",
        127 => "0000000100100111",
        128 => "0000000100101000",
        129 => "0000000100101001",
        130 => "0000000100110000",
        131 => "0000000100110001",
        132 => "0000000100110010",
        133 => "0000000100110011",
        134 => "0000000100110100",
        135 => "0000000100110101",
        136 => "0000000100110110",
        137 => "0000000100110111",
        138 => "0000000100111000",
        139 => "0000000100111001",
        140 => "0000000101000000",
        141 => "0000000101000001",
        142 => "0000000101000010",
        143 => "0000000101000011",
        144 => "0000000101000100",
        145 => "0000000101000101",
        146 => "0000000101000110",
        147 => "0000000101000111",
        148 => "0000000101001000",
        149 => "0000000101001001",
        150 => "0000000101010000",
        151 => "0000000101010001",
        152 => "0000000101010010",
        153 => "0000000101010011",
        154 => "0000000101010100",
        155 => "0000000101010101",
        156 => "0000000101010110",
        157 => "0000000101010111",
        158 => "0000000101011000",
        159 => "0000000101011001",
        160 => "0000000101100000",
        161 => "0000000101100001",
        162 => "0000000101100010",
        163 => "0000000101100011",
        164 => "0000000101100100",
        165 => "0000000101100101",
        166 => "0000000101100110",
        167 => "0000000101100111",
        168 => "0000000101101000",
        169 => "0000000101101001",
        170 => "0000000101110000",
        171 => "0000000101110001",
        172 => "0000000101110010",
        173 => "0000000101110011",
        174 => "0000000101110100",
        175 => "0000000101110101",
        176 => "0000000101110110",
        177 => "0000000101110111",
        178 => "0000000101111000",
        179 => "0000000101111001",
        180 => "0000000110000000",
        181 => "0000000110000001",
        182 => "0000000110000010",
        183 => "0000000110000011",
        184 => "0000000110000100",
        185 => "0000000110000101",
        186 => "0000000110000110",
        187 => "0000000110000111",
        188 => "0000000110001000",
        189 => "0000000110001001",
        190 => "0000000110010000",
        191 => "0000000110010001",
        192 => "0000000110010010",
        193 => "0000000110010011",
        194 => "0000000110010100",
        195 => "0000000110010101",
        196 => "0000000110010110",
        197 => "0000000110010111",
        198 => "0000000110011000",
        199 => "0000000110011001",
        200 => "0000001000000000",
        201 => "0000001000000001",
        202 => "0000001000000010",
        203 => "0000001000000011",
        204 => "0000001000000100",
        205 => "0000001000000101",
        206 => "0000001000000110",
        207 => "0000001000000111",
        208 => "0000001000001000",
        209 => "0000001000001001",
        210 => "0000001000010000",
        211 => "0000001000010001",
        212 => "0000001000010010",
        213 => "0000001000010011",
        214 => "0000001000010100",
        215 => "0000001000010101",
        216 => "0000001000010110",
        217 => "0000001000010111",
        218 => "0000001000011000",
        219 => "0000001000011001",
        220 => "0000001000100000",
        221 => "0000001000100001",
        222 => "0000001000100010",
        223 => "0000001000100011",
        224 => "0000001000100100",
        225 => "0000001000100101",
        226 => "0000001000100110",
        227 => "0000001000100111",
        228 => "0000001000101000",
        229 => "0000001000101001",
        230 => "0000001000110000",
        231 => "0000001000110001",
        232 => "0000001000110010",
        233 => "0000001000110011",
        234 => "0000001000110100",
        235 => "0000001000110101",
        236 => "0000001000110110",
        237 => "0000001000110111",
        238 => "0000001000111000",
        239 => "0000001000111001",
        240 => "0000001001000000",
        241 => "0000001001000001",
        242 => "0000001001000010",
        243 => "0000001001000011",
        244 => "0000001001000100",
        245 => "0000001001000101",
        246 => "0000001001000110",
        247 => "0000001001000111",
        248 => "0000001001001000",
        249 => "0000001001001001",
        250 => "0000001001010000",
        251 => "0000001001010001",
        252 => "0000001001010010",
        253 => "0000001001010011",
        254 => "0000001001010100",
        255 => "0000001001010101"
    );

begin

    process(bin_in)
        variable bcd_out: std_logic_vector(15 downto 0);
    begin
        
        bcd_out := bcd(to_integer(unsigned(bin_in)));

        -- Separar em dígitos BCD
        bcd0 <= bcd_out(3 downto 0);   -- Unidade
        bcd1 <= bcd_out(7 downto 4);   -- Dezena
        bcd2 <= bcd_out(11 downto 8);  -- Centena
        bcd3 <= bcd_out(15 downto 12); -- Milhar
    end process;

end architecture;
